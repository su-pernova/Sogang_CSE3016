`timescale 1ns / 1ps

module buffer(
    input a,
    output y
    );
buf b1(y,a);

endmodule
